blah bolah